/*only takes in clk as an input 
drives itself
get pc next to pc - does the job of pc+4 and mux 
set dummy? 
initialize pcnext as 00000000 feed to pc module 
after pc spits out adress it talks to memory and devides instruction and feeds it */