module testbench(
    
);
endmodule
